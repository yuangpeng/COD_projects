module mccomp(
input			clk,
input			rstn,
input	[4:0]	reg_sel,

output	[31:0]	reg_data
);

	wire	[31:0]	instr;
	wire	[31:0]	PC;
	wire			MemWrite;
	wire	[31:0]	dm_addr;
	wire	[31:0]	dm_din;
	wire	[31:0]	dm_dout;
	
	wire rst = ~rstn;

	// instantiation of single-cycle CPU   
	mccpu U_MCCPU(
		.clk(clk),                 // input:  cpu clock
        .rst(rst),                 // input:  reset
        .instr(instr),             // input:  instruction
        .readdata(dm_dout),        // input:  data to cpu
        .MemWrite(MemWrite),       // output: memory write signal
        .PC(PC),                   // output: PC
        .adr(dm_addr),             // output: address from cpu to memory
        .writedata(dm_din),        // output: data from cpu to memory
        .reg_sel(reg_sel),         // input:  register selection
        .reg_data(reg_data)        // output: register data
    );
         
	// instantiation of data memory  
	dm U_DM(
        .clk(clk),           		// input:  cpu clock
        .DMWr(MemWrite),     		// input:  ram write
        .addr(dm_addr[8:2]), 		// input:  ram address
        .din(dm_din),       		// input:  data to ram
        .dout(dm_dout)      		// output: data from ram
	);
	
endmodule