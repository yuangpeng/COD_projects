`timescale 1ns/1ps

module sll_tb();



endmodule